----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:05:57 02/08/2021 
-- Design Name: 
-- Module Name:    constants - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

package constants is

	type BITMAP1 is array (0 to 88) of std_logic_vector(0 to 339);
	type BITMAP2 is array (0 to 144) of std_logic_vector(0 to 289);
	
	constant logo: BITMAP1 :=
	("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000111111111111111111111111111110000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000000000000000001111",
	"1111100000000000000000000000000000010111111111000000000000000000000000000001111111111111000000000000000000000000000001111111111100000000000000000000000000011111111111111110000000000000000000000000000000000000000001111111111111110000000000000000000000000000011111111111000000000000000000000000000010111111111111111111111111111111111111101111",
	"1111100000000000000000000000000001111111111111100000000000000000000000000001111111111110000000000000000000000000000111111111111110000000000000000000000000000111111111111110000000000000000000000000000000000000000001111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111110000000000000000000000000001111111111100000000000000000000000000000111111111111110000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111110000000000000000000000000001111111111100000000000000000000000000000111111111111110000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111110000000000000000000000000001111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111110000000000000000000000000001111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111110000000000000000000000000001111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111110000000000000000000000000001111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111110000000000000000000000000001111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111110000000000000000000000000001111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111110000000000000000000000000001111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111110000000000000000000000000001111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111110000000000000000000000000001111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111110000000000000000000000000001111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111110000000000000000000000000001111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111100000000000000000000000000001111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000111111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000001111111111111100000000000000000000000000001111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000011111111111110000000000000000000000000000011111111100000000000000000000000000001111111111111111111111111111111111111111111111",
	"1111100000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111110000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111111000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111100000000000000000000000000000111111111111110000000000000000000000000000111111111111110000000000000000000000000000011111111111111000000000000000000000000000000000000000000011111111100000000000000000000000000001111111111111110000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000000000000011111111111100000000000000000000000000000111111111111110000000000000000000000000000011111111111111100000000000000000000000000000000000000000011111111100000000000000000000000000000111111111111100000000000000000000000000001111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111110000000000000000000000000000011111111111111111111111111100000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000001111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111111110000000000000000000000000000011111111111111111111111000000000000000000000000000000000000000000011111111111111111",
	"1111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000111111111111111111111111111110000000000000000000000000000111111111111111111111111100000000000000000000000000000000000000000111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"
	);
	
	constant gOver : BITMAP2 := 
	("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111110000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000000000000011111111110000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000000000000011111111110000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000000000000011111111110000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000000000000011111111110000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000000000000011111111110000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000000000000011111111110000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000000000000011111111110000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000000000000011111111110000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000000000000011111111110000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000011111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111110000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111110000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111110000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111110000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111110000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111110000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111110000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111110000000000000000000000000000111111111000000000000000000111111111111111111111111111100000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000001111111100000000001111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000001111111100000000011111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000001111111100000000011111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000001111111100000000011111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000001111111100000000011111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000001111111100000000011111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000001111111100000000011111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000001111111100000000011111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000001111111100000000011111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000011111111100000000000000000001111111110000000011111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111100000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000001111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000111111111111111111111111111111111111111111111111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111110000000000000000000000000000000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111100000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11111111111100000000000000000000000000000000000000000000001111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000111111111111",
	"11101001001100000000001111111111111111111111111110000000000100000001111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111000000000010000010111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111100000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111100000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111100000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111100000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111100000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111100000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111100000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111100000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111100000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111100000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111100000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111000000000000000000111111111111111111111111111000000000000000000011111111100000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111000000000011111111111111111101111111000000000011111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111000000000011111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111000000000000000000111111111100000000000000000011111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000000000000011111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111000000000000000000000000000111111111111",
	"11100000000000000000001111111111111111111111111110000000000000000000111111111111111111111111111000000000000000000000000000111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000111111111000000000000000000000000000111111111111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11111111111110000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000111111111111111111000000000000000000000000000111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
	"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"
	);
end constants;

